module full_sub_tb;

reg A, B, Bin;
wire D, Bout;

full_sub uut (
    .A(A),
    .B(B),
    .Bin(Bin),
    .D(D),
    .Bout(Bout)
);

initial begin
    $dumpfile("full_sub_tb.vcd");
    $dumpvars(0, full_sub_tb);
end

initial begin
    A=0; B=0; Bin=0;
    #10 A=0; B=0; Bin=1;
    #10 A=0; B=1; Bin=0;
    #10 A=0; B=1; Bin=1;
    #10 A=1; B=0; Bin=0;
    #10 A=1; B=0; Bin=1;
    #10 A=1; B=1; Bin=0;
    #10 A=1; B=1; Bin=1;
    #10 $finish;
end

endmodule


